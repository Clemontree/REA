05 21 2021 10 51 04     1     0    48    53    51     2     7     3   114.7   188.4   188.9   303.2   155.9   114.7   188.4   188.9   303.2   155.9
05 21 2021 11 21 33     2     0    47    48    50     5     4     3   186.6   185.6   130.4   300.0   152.7   186.6   185.6   130.4   300.3   152.8
05 21 2021 13 45 53     3     0    47    50    51     2     4     3   126.8   170.0   178.5     0.0     0.0   126.8   170.0   178.5     0.0     0.0
