05 20 2021 15 14 26     1     0    48    51    51     1     2     4   208.8   192.3   191.2   307.9   160.7   208.8   192.3   191.2   307.9   160.7
