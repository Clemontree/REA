06 05 2021 13 10 58     1     0    52    53    57     7     1     4   147.7   168.6   166.7   272.0   123.3   147.7   168.6   166.7   271.5   123.1
06 05 2021 13 27 58     2     0    47    47    50     2     3     6   147.5   167.3   164.9     0.0     0.0   147.5   167.3   164.9     0.0     0.0
06 05 2021 14 07 00     3     0    45    46    45     1     5     8    -1.0   115.2    -1.0     0.0     0.0    -1.0   115.2    -1.0     0.0     0.0
