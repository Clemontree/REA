06 05 2021 14 42 03     1     0    45    45    45     2     5     7   114.5   111.4   112.7   184.4    35.3   114.5   111.4   112.7   184.4    35.3
