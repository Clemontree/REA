10 15 2020 08 47 22     1     0    45    47    47     1     4     4   188.5   183.1   186.8   300.6   153.8   188.5   183.1   186.8   300.6   153.8
10 15 2020 08 48 23     2     0    45    46    47     7     8     3   188.2   183.5   119.3     0.0     0.0   188.2   183.5   119.3     0.0     0.0
10 15 2020 09 58 43     3     0    45    47    47     3     5     7   177.9   176.0   178.6   284.7   137.9   177.9   176.0   178.6   284.7   137.9
10 15 2020 10 45 14     4     0    46    49    49     4     6     1   177.0   171.6   178.4   284.7   137.9   177.0   171.6   178.4   284.7   137.9
10 15 2020 10 49 02     5     0    45    47    47     6     3     3   177.3   189.1   112.9     0.0     0.0   177.3   189.1   112.9     0.0     0.0
10 15 2020 10 56 32     6     0    45    46    47     5     1     8   176.7   178.9   182.8     0.0     0.0   176.7   178.9   182.8     0.0     0.0
