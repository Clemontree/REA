04 29 2021 10 38 39     1     0    50    50    53     5     5     3   253.4   217.7   218.4   348.2   202.1   253.4   217.7   218.4   348.2   202.1
