05 21 2021 14 28 58     1     0    46    48    49     3     3     6   117.8   111.1   113.3     0.0     0.0   117.8   111.1   113.3     0.0     0.0
