06 05 2021 15 45 36     1     0    46    46    47     4     6    12   119.3   117.8   106.8   192.5    43.5   119.3   117.8   106.8   192.5    43.5
