04 21 2021 11 31 09     1     0    45    46    47     7     1     3   239.4   249.3   237.9   384.9   236.7   239.4   249.3   237.9   384.9   236.7
