04 29 2021 09 53 37     1     0    50    50    53     6     8     7   252.6   227.8   230.4     0.0     0.0   252.6   227.8   230.4     0.0     0.0
